// Code your design here
`include "platform.sv"
`include "definitions.sv"
`include "alu.sv"
`include "cpu.sv"
`include "top.sv"
`include "ram_sim.v"
`include "rom_sim.v"
